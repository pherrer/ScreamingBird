--WORK IN PROGRESS
